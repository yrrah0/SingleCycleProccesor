library verilog;
use verilog.vl_types.all;
entity enARdFF_1_vlg_vec_tst is
end enARdFF_1_vlg_vec_tst;
