library verilog;
use verilog.vl_types.all;
entity ProcessorMIPSBenchTest_vlg_vec_tst is
end ProcessorMIPSBenchTest_vlg_vec_tst;
