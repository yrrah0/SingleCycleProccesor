library verilog;
use verilog.vl_types.all;
entity fullAdder32bit_vlg_vec_tst is
end fullAdder32bit_vlg_vec_tst;
