library verilog;
use verilog.vl_types.all;
entity ProcessorControl_vlg_vec_tst is
end ProcessorControl_vlg_vec_tst;
