library verilog;
use verilog.vl_types.all;
entity TopLevelMIPS_vlg_vec_tst is
end TopLevelMIPS_vlg_vec_tst;
