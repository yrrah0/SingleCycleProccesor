library verilog;
use verilog.vl_types.all;
entity PCAddTest_vlg_vec_tst is
end PCAddTest_vlg_vec_tst;
