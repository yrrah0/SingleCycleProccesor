library verilog;
use verilog.vl_types.all;
entity ALUControl_vlg_vec_tst is
end ALUControl_vlg_vec_tst;
