library verilog;
use verilog.vl_types.all;
entity CompTest_vlg_vec_tst is
end CompTest_vlg_vec_tst;
