library verilog;
use verilog.vl_types.all;
entity testBlockFile_vlg_vec_tst is
end testBlockFile_vlg_vec_tst;
