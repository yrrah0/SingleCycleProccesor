library verilog;
use verilog.vl_types.all;
entity testBlock_vlg_vec_tst is
end testBlock_vlg_vec_tst;
