library verilog;
use verilog.vl_types.all;
entity testBlockUnit_vlg_vec_tst is
end testBlockUnit_vlg_vec_tst;
