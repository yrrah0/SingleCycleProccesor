library verilog;
use verilog.vl_types.all;
entity instructionPCTest_vlg_vec_tst is
end instructionPCTest_vlg_vec_tst;
